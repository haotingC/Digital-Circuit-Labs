module t_Lab2_decoder_5x32;
      wire   [31:0]Dout;
      reg    [4:0]A;
      reg    enable;

      Lab2_decoder_5x32    d1(Dout, A, enable);
      

      initial begin 
              A[4]=1'b0; A[3]=1'b0; A[2]=1'b0; A[1]=1'b0; A[0]=1'b0; enable=1'b0;
              #100 A[4]=1'b0; A[3]=1'b0; A[2]=1'b0; A[1]=1'b0; A[0]=1'b1; enable=1'b0;
              #100 A[4]=1'b0; A[3]=1'b0; A[2]=1'b0; A[1]=1'b1; A[0]=1'b0; enable=1'b0;
              #100 A[4]=1'b0; A[3]=1'b0; A[2]=1'b0; A[1]=1'b1; A[0]=1'b1; enable=1'b0;
              #100 A[4]=1'b0; A[3]=1'b0; A[2]=1'b1; A[1]=1'b0; A[0]=1'b0; enable=1'b0;
              #100 A[4]=1'b0; A[3]=1'b0; A[2]=1'b1; A[1]=1'b0; A[0]=1'b1; enable=1'b0;
              #100 A[4]=1'b0; A[3]=1'b0; A[2]=1'b1; A[1]=1'b1; A[0]=1'b0; enable=1'b0;
              #100 A[4]=1'b0; A[3]=1'b0; A[2]=1'b1; A[1]=1'b1; A[0]=1'b1; enable=1'b0;
              #100 A[4]=1'b0; A[3]=1'b1; A[2]=1'b0; A[1]=1'b0; A[0]=1'b0; enable=1'b0;
              #100 A[4]=1'b0; A[3]=1'b1; A[2]=1'b0; A[1]=1'b0; A[0]=1'b1; enable=1'b0;
              #100 A[4]=1'b0; A[3]=1'b1; A[2]=1'b0; A[1]=1'b1; A[0]=1'b0; enable=1'b0;
              #100 A[4]=1'b0; A[3]=1'b1; A[2]=1'b0; A[1]=1'b1; A[0]=1'b1; enable=1'b0;
              #100 A[4]=1'b0; A[3]=1'b1; A[2]=1'b1; A[1]=1'b0; A[0]=1'b0; enable=1'b0;
              #100 A[4]=1'b0; A[3]=1'b1; A[2]=1'b1; A[1]=1'b0; A[0]=1'b1; enable=1'b0;
              #100 A[4]=1'b0; A[3]=1'b1; A[2]=1'b1; A[1]=1'b1; A[0]=1'b0; enable=1'b0;
              #100 A[4]=1'b0; A[3]=1'b1; A[2]=1'b1; A[1]=1'b1; A[0]=1'b1; enable=1'b0;
              #100 A[4]=1'b1; A[3]=1'b0; A[2]=1'b0; A[1]=1'b0; A[0]=1'b0; enable=1'b0;
              #100 A[4]=1'b1; A[3]=1'b0; A[2]=1'b0; A[1]=1'b0; A[0]=1'b1; enable=1'b0;
              #100 A[4]=1'b1; A[3]=1'b0; A[2]=1'b0; A[1]=1'b1; A[0]=1'b0; enable=1'b0;
              #100 A[4]=1'b1; A[3]=1'b0; A[2]=1'b0; A[1]=1'b1; A[0]=1'b1; enable=1'b0;
              #100 A[4]=1'b1; A[3]=1'b0; A[2]=1'b1; A[1]=1'b0; A[0]=1'b0; enable=1'b0;
              #100 A[4]=1'b1; A[3]=1'b0; A[2]=1'b1; A[1]=1'b0; A[0]=1'b1; enable=1'b0;
              #100 A[4]=1'b1; A[3]=1'b0; A[2]=1'b1; A[1]=1'b1; A[0]=1'b0; enable=1'b0;
              #100 A[4]=1'b1; A[3]=1'b0; A[2]=1'b1; A[1]=1'b1; A[0]=1'b1; enable=1'b0;
              #100 A[4]=1'b1; A[3]=1'b1; A[2]=1'b0; A[1]=1'b0; A[0]=1'b0; enable=1'b0;
              #100 A[4]=1'b1; A[3]=1'b1; A[2]=1'b0; A[1]=1'b0; A[0]=1'b1; enable=1'b0;
              #100 A[4]=1'b1; A[3]=1'b1; A[2]=1'b0; A[1]=1'b1; A[0]=1'b0; enable=1'b0;
              #100 A[4]=1'b1; A[3]=1'b1; A[2]=1'b0; A[1]=1'b1; A[0]=1'b1; enable=1'b0;
              #100 A[4]=1'b1; A[3]=1'b1; A[2]=1'b1; A[1]=1'b0; A[0]=1'b0; enable=1'b0;
              #100 A[4]=1'b1; A[3]=1'b1; A[2]=1'b1; A[1]=1'b0; A[0]=1'b1; enable=1'b0;
              #100 A[4]=1'b1; A[3]=1'b1; A[2]=1'b1; A[1]=1'b1; A[0]=1'b0; enable=1'b0;
              #100 A[4]=1'b1; A[3]=1'b1; A[2]=1'b1; A[1]=1'b1; A[0]=1'b1; enable=1'b0;

              #100 A[4]=1'b0; A[3]=1'b0; A[2]=1'b0; A[1]=1'b0; A[0]=1'b0; enable=1'b1;
              #100 A[4]=1'b0; A[3]=1'b0; A[2]=1'b0; A[1]=1'b0; A[0]=1'b1; enable=1'b1;
              #100 A[4]=1'b0; A[3]=1'b0; A[2]=1'b0; A[1]=1'b1; A[0]=1'b0; enable=1'b1;
              #100 A[4]=1'b0; A[3]=1'b0; A[2]=1'b0; A[1]=1'b1; A[0]=1'b1; enable=1'b1;
              #100 A[4]=1'b0; A[3]=1'b0; A[2]=1'b1; A[1]=1'b0; A[0]=1'b0; enable=1'b1;
              #100 A[4]=1'b0; A[3]=1'b0; A[2]=1'b1; A[1]=1'b0; A[0]=1'b1; enable=1'b1;
              #100 A[4]=1'b0; A[3]=1'b0; A[2]=1'b1; A[1]=1'b1; A[0]=1'b0; enable=1'b1;
              #100 A[4]=1'b0; A[3]=1'b0; A[2]=1'b1; A[1]=1'b1; A[0]=1'b1; enable=1'b1;
              #100 A[4]=1'b0; A[3]=1'b1; A[2]=1'b0; A[1]=1'b0; A[0]=1'b0; enable=1'b1;
              #100 A[4]=1'b0; A[3]=1'b1; A[2]=1'b0; A[1]=1'b0; A[0]=1'b1; enable=1'b1;
              #100 A[4]=1'b0; A[3]=1'b1; A[2]=1'b0; A[1]=1'b1; A[0]=1'b0; enable=1'b1;
              #100 A[4]=1'b0; A[3]=1'b1; A[2]=1'b0; A[1]=1'b1; A[0]=1'b1; enable=1'b1;
              #100 A[4]=1'b0; A[3]=1'b1; A[2]=1'b1; A[1]=1'b0; A[0]=1'b0; enable=1'b1;
              #100 A[4]=1'b0; A[3]=1'b1; A[2]=1'b1; A[1]=1'b0; A[0]=1'b1; enable=1'b1;
              #100 A[4]=1'b0; A[3]=1'b1; A[2]=1'b1; A[1]=1'b1; A[0]=1'b0; enable=1'b1;
              #100 A[4]=1'b0; A[3]=1'b1; A[2]=1'b1; A[1]=1'b1; A[0]=1'b1; enable=1'b1;
              #100 A[4]=1'b1; A[3]=1'b0; A[2]=1'b0; A[1]=1'b0; A[0]=1'b0; enable=1'b1;
              #100 A[4]=1'b1; A[3]=1'b0; A[2]=1'b0; A[1]=1'b0; A[0]=1'b1; enable=1'b1;
              #100 A[4]=1'b1; A[3]=1'b0; A[2]=1'b0; A[1]=1'b1; A[0]=1'b0; enable=1'b1;
              #100 A[4]=1'b1; A[3]=1'b0; A[2]=1'b0; A[1]=1'b1; A[0]=1'b1; enable=1'b1;
              #100 A[4]=1'b1; A[3]=1'b0; A[2]=1'b1; A[1]=1'b0; A[0]=1'b0; enable=1'b1;
              #100 A[4]=1'b1; A[3]=1'b0; A[2]=1'b1; A[1]=1'b0; A[0]=1'b1; enable=1'b1;
              #100 A[4]=1'b1; A[3]=1'b0; A[2]=1'b1; A[1]=1'b1; A[0]=1'b0; enable=1'b1;
              #100 A[4]=1'b1; A[3]=1'b0; A[2]=1'b1; A[1]=1'b1; A[0]=1'b1; enable=1'b1;
              #100 A[4]=1'b1; A[3]=1'b1; A[2]=1'b0; A[1]=1'b0; A[0]=1'b0; enable=1'b1;
              #100 A[4]=1'b1; A[3]=1'b1; A[2]=1'b0; A[1]=1'b0; A[0]=1'b1; enable=1'b1;
              #100 A[4]=1'b1; A[3]=1'b1; A[2]=1'b0; A[1]=1'b1; A[0]=1'b0; enable=1'b1;
              #100 A[4]=1'b1; A[3]=1'b1; A[2]=1'b0; A[1]=1'b1; A[0]=1'b1; enable=1'b1;
              #100 A[4]=1'b1; A[3]=1'b1; A[2]=1'b1; A[1]=1'b0; A[0]=1'b0; enable=1'b1;
              #100 A[4]=1'b1; A[3]=1'b1; A[2]=1'b1; A[1]=1'b0; A[0]=1'b1; enable=1'b1;
              #100 A[4]=1'b1; A[3]=1'b1; A[2]=1'b1; A[1]=1'b1; A[0]=1'b0; enable=1'b1;
              #100 A[4]=1'b1; A[3]=1'b1; A[2]=1'b1; A[1]=1'b1; A[0]=1'b1; enable=1'b1;
      end 
      initial #6400 $finish;
endmodule 
